* Netlista sumatora
.subckt SUMATOR A B C SUM CARRY VDD VSS


********************Blok CARRY
*Tablica PMOS
M1 s1 A VDD VDD PCH L=0.065u W=0.94u M=1
M2 s1 B VDD VDD PCH L=0.065u W=0.94u M=1
M3 s2 B s1 VDD PCH L=0.065u W=0.94u M=1
M4 Ca C s1 VDD PCH L=0.065u W=0.94u M=1
M5 Ca A s2 VDD PCH L=0.065u W=0.94u M=1

*Tablica NMOS
M6 s1 A VDD VDD NCH L=0.065u W=0.2u M=1
M7 s1 B VDD VDD NCH L=0.065u W=0.2u M=1
M8 s2 B s1 VDD NCH L=0.065u W=0.2u M=1
M9 Ca C s1 VDD NCH L=0.065u W=0.2u M=1
M10 Ca A s2 VDD NCH L=0.065u W=0.2u M=1

*INV
*M11 s1 A VDD VDD PCH L=0.065u W=0.94u M=1
*M12 s1 A VDD VDD PCH L=0.065u W=0.94u M=1
...

********************BLOK SUM
*Tablica PMOS
M13 s5 A VDD VDD PCH L=0.065u W=0.94u M=1
M14 s5 B VDD VDD PCH L=0.065u W=0.94u M=1
M15 s5 C VDD VDD PCH L=0.065u W=0.94u M=1
M16 s6 A s5 VDD PCH L=0.065u W=0.94u M=1
M17 s7 B s6 VDD PCH L=0.065u W=0.94u M=1
M18 S C s7 VDD PCH L=0.065u W=0.94u M=1
M19 S Ca s5 VDD PCH L=0.065u W=0.94u M=1

*Tablica NMOS
M20 s1 A VDD VDD NCH L=0.065u W=0.2u M=1
M21 s1 B VDD VDD NCH L=0.065u W=0.2u M=1
M22 s2 B s1 VDD NCH L=0.065u W=0.2u M=1
M23 Ca C s1 VDD NCH L=0.065u W=0.2u M=1
M24 Ca A s2 VDD NCH L=0.065u W=0.2u M=1
M25 s1 A VDD VDD NCH L=0.065u W=0.2u M=1
M26 s1 B VDD VDD NCH L=0.065u W=0.2u M=1


*INV
M27 s1 A VDD VDD PCH L=0.065u W=0.94u M=1
M28 s1 B VDD VDD PCH L=0.065u W=0.94u M=1


.ends