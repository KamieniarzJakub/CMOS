.include sumator.sp

.subckt 4BITOWY A1 A2 A3 A4 B1 B2 B3 B4 Cin S1 S2 S3 S4 Cout VDD VSS
XSUM1 A1 B1 Cin S1 C2 VDD VSS SUMATOR
XSUM2 A2 B2 C2 S2 C3 VDD VSS SUMATOR
XSUM3 A3 B3 C3 S3 C4 VDD VSS SUMATOR
XSUM4 A4 B4 C4 S4 Cout VDD VSS SUMATOR
.ends
